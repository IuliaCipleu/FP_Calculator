package CONSTANTS is
	constant NumBit : integer := 24;	
	
end package CONSTANTS;